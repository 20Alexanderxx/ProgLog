--Verhaltensmodell 
library ieee; 
use ieee.std_logic_1164.all; 

entity siebenseg is 
port( b : in std_logic_vector(3 downto 0); -- b3 to b0 
    ltn, bin : in std_logic; 
    hex : out std_logic_vector(0 to 6)); -- hex00..hex06 
end siebenseg; 
 
 architecture behavior of siebenseg is 
 begin 
 
    pl: process ( ltn, bin, b ) 
    begin 
        if ( ltn = '1' and bin = '0' ) then 
            case b is 
                --segmente abcdefg 
                when "0000"=> hex <="0000001"; -- 0 
                when "0001"=> hex <="1001111"; -- 1 
                when "0010"=> hex <="0010010"; -- 2 
                when "0011"=> hex <="0000110"; -- 3 
                when "0100"=> hex <="1001100"; -- 4 
                when "0101"=> hex <="0100100"; -- 5 
                when "0110"=> hex <="0100000"; -- 6 
                when "0111"=> hex <="0001111"; -- 7 
                when "1000"=> hex <="0000000"; -- 8 
                when "1001"=> hex <="0000100"; -- 9 
                when "1010"=> hex <="0001000"; -- A -> 10 
                when "1011"=> hex <="1100000"; -- b -> 11 
                when "1100"=> hex <="0110001"; -- C -> 12 
                when "1101"=> hex <="1000010"; -- d -> 13 
                when "1110"=> hex <="0110000"; -- E -> 14 
                when "1111"=> hex <="0111000"; -- F -> 15 
                when others=> hex <="0000000"; -- should not 
            end case; 
        elsif ( ltn = '0' and bin = '1' ) then 
            hex <= "0000000"; 
        elsif ( ltn = '0' and bin = '0' ) then 
            hex <= "1111111"; 
        else 
            -- dummy 
            hex <= "1111111"; 
        end if; 
    end process pl; 
 
 end behavior; 