Library ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity bcd_tb is
end bcd_tb;

architecture testbench of bcd_tb is
component bcd 
	port(	b : in std_logic_vector(3 downto 0);
			ltn, bin : in std_logic; 
			hex : out std_logic_vector(0 to 6));
end component;

signal b_s : std_logic_vector(3 downto 0);
signal ltn_s, bin_s : std_logic;
signal hex_s : std_logic_vector(0 to 6);

begin
dut: bcd
port map (b_s, ltn_s, bin_s, hex_s);
process
begin
	ltn_s <= '0'; bin_s <= '0'; b_s <= "0000";
	wait for 1ns;
	b_s <= "0001";
	wait for 1ns;
	b_s <= "0010";
	wait for 1ns;
	b_s <= "0011";
	wait for 1ns;
	b_s <= "0100";
	wait for 1ns;
	b_s <= "0101";
	wait for 1ns;
	b_s <= "0110";
	wait for 1ns;
	b_s <= "0111";
	wait for 1ns;
	b_s <= "1000";
	wait for 1ns;
	b_s <= "1001";
	wait for 1ns;
	b_s <= "1010";
	wait for 1ns;
	b_s <= "1011";
	wait for 1ns;
	b_s <= "1100";
	wait for 1ns;
	b_s <= "1101";
	wait for 1ns;
	b_s <= "1110";
	wait for 1ns;
	b_s <= "1111";
	wait for 1ns;
	ltn_s <= '0'; bin_s <= '1'; b_s <= "0000";
	wait for 1ns;
	b_s <= "0001";
	wait for 1ns;
	b_s <= "0010";
	wait for 1ns;
	b_s <= "0011";
	wait for 1ns;
	b_s <= "0100";
	wait for 1ns;
	b_s <= "0101";
	wait for 1ns;
	b_s <= "0110";
	wait for 1ns;
	b_s <= "0111";
	wait for 1ns;
	b_s <= "1000";
	wait for 1ns;
	b_s <= "1001";
	wait for 1ns;
	b_s <= "1010";
	wait for 1ns;
	b_s <= "1011";
	wait for 1ns;
	b_s <= "1100";
	wait for 1ns;
	b_s <= "1101";
	wait for 1ns;
	b_s <= "1110";
	wait for 1ns;
	b_s <= "1111";
	wait for 1ns;
	ltn_s <= '1'; bin_s <= '0'; b_s <= "0000";
	wait for 1ns;
	b_s <= "0001";
	wait for 1ns;
	b_s <= "0010";
	wait for 1ns;
	b_s <= "0011";
	wait for 1ns;
	b_s <= "0100";
	wait for 1ns;
	b_s <= "0101";
	wait for 1ns;
	b_s <= "0110";
	wait for 1ns;
	b_s <= "0111";
	wait for 1ns;
	b_s <= "1000";
	wait for 1ns;
	b_s <= "1001";
	wait for 1ns;
	b_s <= "1010";
	wait for 1ns;
	b_s <= "1011";
	wait for 1ns;
	b_s <= "1100";
	wait for 1ns;
	b_s <= "1101";
	wait for 1ns;
	b_s <= "1110";
	wait for 1ns;
	b_s <= "1111";
	wait for 1ns;
	ltn_s <= '1'; bin_s <= '1'; b_s <= "0000";
	wait for 1ns;
	b_s <= "0001";
	wait for 1ns;
	b_s <= "0010";
	wait for 1ns;
	b_s <= "0011";
	wait for 1ns;
	b_s <= "0100";
	wait for 1ns;
	b_s <= "0101";
	wait for 1ns;
	b_s <= "0110";
	wait for 1ns;
	b_s <= "0111";
	wait for 1ns;
	b_s <= "1000";
	wait for 1ns;
	b_s <= "1001";
	wait for 1ns;
	b_s <= "1010";
	wait for 1ns;
	b_s <= "1011";
	wait for 1ns;
	b_s <= "1100";
	wait for 1ns;
	b_s <= "1101";
	wait for 1ns;
	b_s <= "1110";
	wait for 1ns;
	b_s <= "1111";
	wait for 1ns;
	wait;
end process;
end testbench;